
-- Code your design here
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith
ENTITY FA1 is 
	port(a,b,ci:in std_logic;s,cout:out std_logic);
end FA1;
architecture structural of FA1 is

begin
end structural; 