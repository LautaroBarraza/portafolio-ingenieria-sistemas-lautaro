library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity Registers is
	Generic (
		B: integer := 32; -- numero de bits del registro
		W: integer := 5  -- numero de bits de direcciones
	);
	Port(reg1_rd  : in std_logic_vector(W-1 downto 0);
		 reg2_rd  : in std_logic_vector(W-1 downto 0);
		 reg_wr   : in std_logic_vector(W-1 downto 0);
		 data_wr  : in std_logic_vector(B-1 downto 0);
		 wr       : in std_logic;
		 reset    : in std_logic;
		 clk      : in std_logic;
		 data1_rd : out std_logic_vector(B-1 downto 0);
		 data2_rd : out std_logic_vector(B-1 downto 0)
);
end Registers;

architecture PRACTICA of Registers is
	type reg_file_type is array(0 to (2**W)-1) of std_logic_vector(B-1 downto 0);
	signal reg_outputs: reg_file_type:= (others => (others => '0')); 
	
begin
	data1_rd <= reg_outputs(conv_integer(reg1_rd)) when reg1_rd /= x"00000000" else x"00000000";
	data2_rd <= reg_outputs(conv_integer(reg2_rd)) when reg2_rd /= x"00000000" else x"00000000";
    
	writting:process(clk,reset)
    begin
        if reset='1' then
          	reg_outputs <= (others => (others => '0'));
        elsif falling_edge(clk) then
        	if(wr='1') then
            	reg_outputs(conv_integer(reg_wr)) <= data_wr;
          	end if;
      	end if;
    end process; 
end PRACTICA;
